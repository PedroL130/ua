library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity NoisyTriangSignal_ROM_256x8 is
   port(address : in  std_logic_vector(7 downto 0);
        dataOut : out std_logic_vector(7 downto 0));
end NoisyTriangSignal_ROM_256x8;

architecture Behavioral of NoisyTriangSignal_ROM_256x8 is
   subtype TDataWord is std_logic_vector(7 downto 0);
   type TROM is array (0 to 255) of TDataWord;
	-- Input Signal ROM
   constant c_memory: TROM := (
	"11000000",
	"11000010",
	"11000100",
	"11000110",
	"11001001",
	"11001011",
	"11001101",
	"11001111",
	"11011101",
	"11010011",
	"11010101",
	"11010111",
	"11011010",
	"11011100",
	"11011110",
	"11100000",
	"11100010",
	"11100100",
	"11100110",
	"11101001",
	"11101011",
	"11101101",
	"11101111",
	"11110001",
	"11110011",
	"11110101",
	"11110111",
	"11111000",
	"11111100",
	"11111110",
	"00000000",
	"00000010",
	"00000011",
	"00000110",
	"00001001",
	"00001011",
	"00001101",
	"00010011",
	"00010001",
	"00010011",
	"00010101",
	"00010111",
	"00100000",
	"00011100",
	"00100101",
	"00100000",
	"00011010",
	"00100100",
	"00100110",
	"00101001",
	"00101011",
	"00101101",
	"00100011",
	"00110001",
	"00110011",
	"00110101",
	"00110111",
	"01001000",
	"00111100",
	"01001101",
	"01000000",
	"00111110",
	"00111100",
	"00111010",
	"00110111",
	"00101000",
	"00110011",
	"00110001",
	"00101111",
	"00101101",
	"00101011",
	"00101001",
	"00100110",
	"00100100",
	"00100010",
	"00101000",
	"00011110",
	"00011100",
	"00011010",
	"00010111",
	"00010101",
	"00010011",
	"00010001",
	"00001111",
	"00001101",
	"00001011",
	"00001001",
	"00000110",
	"00000101",
	"00000010",
	"00000000",
	"11111110",
	"11111100",
	"11111010",
	"11110111",
	"11110101",
	"11110011",
	"11110001",
	"11101111",
	"11101101",
	"11100101",
	"11101001",
	"11100110",
	"11100100",
	"11100010",
	"11100000",
	"11011110",
	"11011100",
	"11011010",
	"11010111",
	"11010101",
	"11011110",
	"11000101",
	"11001111",
	"11001101",
	"11001011",
	"11001001",
	"11000110",
	"11000100",
	"11000010",
	"11000000",
	"11000010",
	"11000100",
	"11000110",
	"11001001",
	"11001011",
	"11001101",
	"11011011",
	"11010001",
	"11010011",
	"11010101",
	"11010111",
	"11100011",
	"11011100",
	"11011110",
	"11100000",
	"11011011",
	"11100100",
	"11101101",
	"11101001",
	"11101011",
	"11101101",
	"11101111",
	"11110001",
	"11110011",
	"11110101",
	"11110111",
	"11111010",
	"11111100",
	"11111110",
	"00000000",
	"00000010",
	"00000101",
	"00000110",
	"00001001",
	"00001011",
	"00001101",
	"00001111",
	"00010001",
	"00010011",
	"00010101",
	"00010010",
	"00011010",
	"00010101",
	"00011110",
	"00100000",
	"00100010",
	"00011011",
	"00100110",
	"00011110",
	"00101011",
	"00101101",
	"00101111",
	"00110001",
	"00110011",
	"00110101",
	"01000101",
	"00111010",
	"00111100",
	"00101110",
	"01000000",
	"00111110",
	"00111100",
	"01001000",
	"00110111",
	"00110101",
	"00110011",
	"00110001",
	"00101111",
	"00101101",
	"00101011",
	"00101001",
	"00100110",
	"00100100",
	"00100010",
	"00100000",
	"00011110",
	"00011100",
	"00011010",
	"00010111",
	"00010101",
	"00010011",
	"00010001",
	"00001011",
	"00001101",
	"00001011",
	"00001001",
	"00000110",
	"00000100",
	"00000010",
	"00000000",
	"11111110",
	"11111100",
	"11111010",
	"11110111",
	"11110101",
	"11110110",
	"11110001",
	"11110011",
	"11101101",
	"11101011",
	"11101001",
	"11100110",
	"11100100",
	"11100010",
	"11100000",
	"11011110",
	"11011100",
	"11011010",
	"11010111",
	"11010101",
	"11010011",
	"11010001",
	"11001111",
	"11001101",
	"10111101",
	"11001001",
	"11000110",
	"11000100",
	"10110011",
	"11000000",
	"11000010",
	"11000100",
	"11000110",
	"11001001",
	"10111101",
	"11001101",
	"11001111",
	"11000101",
	"11010011",
	"11100000",
	"11010111",
	"11011010",
	"11010011",
	"11011110",
	"11100000"
	);

begin
   dataOut <= c_memory(to_integer(unsigned(address)));
end Behavioral;
